//
// Created by Kumonda221 (Ding Haonan) on 2024/03/20
//

`define         PutFullData         0
`define         PutPartialData      1
`define         ArithmeticData      2
`define         LogicalData         3
`define         Get                 4
`define         Intent              5
`define         AcquireBlock        6
`define         AcquirePerm         7

`define         ProbeBlock          6
`define         ProbePerm           7

`define         AccessAck           0
`define         AccessAckData       1
`define         HintAck             2
`define         ProbeAck            4
`define         ProbeAckData        5
`define         Release             6
`define         ReleaseData         7

`define         Grant               4
`define         GrantData           5
`define         ReleaseAck          6

`define         GrantAck            0
