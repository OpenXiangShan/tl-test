`timescale 1ns/1ps

module tb_top(
  input wire clock,
  input wire reset
);
  `include "tb_signals.v"

  assign io_clock = clock;
  assign io_reset = reset;
  XSTop l_soc(
    .s_dma_aw_ready(s_dma_aw_ready),
    .s_dma_aw_valid(s_dma_aw_valid),
    .s_dma_aw_id(s_dma_aw_id),
    .s_dma_aw_addr(s_dma_aw_addr),
    .s_dma_aw_len(s_dma_aw_len),
    .s_dma_aw_size(s_dma_aw_size),
    .s_dma_aw_burst(s_dma_aw_burst),
    .s_dma_aw_lock(s_dma_aw_lock),
    .s_dma_aw_cache(s_dma_aw_cache),
    .s_dma_aw_prot(s_dma_aw_prot),
    .s_dma_aw_qos(s_dma_aw_qos),
    .s_dma_w_ready(s_dma_w_ready),
    .s_dma_w_valid(s_dma_w_valid),
    .s_dma_w_data(s_dma_w_data),
    .s_dma_w_strb(s_dma_w_strb),
    .s_dma_w_last(s_dma_w_last),
    .s_dma_b_ready(s_dma_b_ready),
    .s_dma_b_valid(s_dma_b_valid),
    .s_dma_b_id(s_dma_b_id),
    .s_dma_b_resp(s_dma_b_resp),
    .s_dma_ar_ready(s_dma_ar_ready),
    .s_dma_ar_valid(s_dma_ar_valid),
    .s_dma_ar_id(s_dma_ar_id),
    .s_dma_ar_addr(s_dma_ar_addr),
    .s_dma_ar_len(s_dma_ar_len),
    .s_dma_ar_size(s_dma_ar_size),
    .s_dma_ar_burst(s_dma_ar_burst),
    .s_dma_ar_lock(s_dma_ar_lock),
    .s_dma_ar_cache(s_dma_ar_cache),
    .s_dma_ar_prot(s_dma_ar_prot),
    .s_dma_ar_qos(s_dma_ar_qos),
    .s_dma_r_ready(s_dma_r_ready),
    .s_dma_r_valid(s_dma_r_valid),
    .s_dma_r_id(s_dma_r_id),
    .s_dma_r_data(s_dma_r_data),
    .s_dma_r_resp(s_dma_r_resp),
    .s_dma_r_last(s_dma_r_last),
    .m_peripheral_aw_ready(m_peripheral_aw_ready),
    .m_peripheral_aw_valid(m_peripheral_aw_valid),
    .m_peripheral_aw_id(m_peripheral_aw_id),
    .m_peripheral_aw_addr(m_peripheral_aw_addr),
    .m_peripheral_aw_len(m_peripheral_aw_len),
    .m_peripheral_aw_size(m_peripheral_aw_size),
    .m_peripheral_aw_burst(m_peripheral_aw_burst),
    .m_peripheral_aw_lock(m_peripheral_aw_lock),
    .m_peripheral_aw_cache(m_peripheral_aw_cache),
    .m_peripheral_aw_prot(m_peripheral_aw_prot),
    .m_peripheral_aw_qos(m_peripheral_aw_qos),
    .m_peripheral_w_ready(m_peripheral_w_ready),
    .m_peripheral_w_valid(m_peripheral_w_valid),
    .m_peripheral_w_data(m_peripheral_w_data),
    .m_peripheral_w_strb(m_peripheral_w_strb),
    .m_peripheral_w_last(m_peripheral_w_last),
    .m_peripheral_b_ready(m_peripheral_b_ready),
    .m_peripheral_b_valid(m_peripheral_b_valid),
    .m_peripheral_b_id(m_peripheral_b_id),
    .m_peripheral_b_resp(m_peripheral_b_resp),
    .m_peripheral_ar_ready(m_peripheral_ar_ready),
    .m_peripheral_ar_valid(m_peripheral_ar_valid),
    .m_peripheral_ar_id(m_peripheral_ar_id),
    .m_peripheral_ar_addr(m_peripheral_ar_addr),
    .m_peripheral_ar_len(m_peripheral_ar_len),
    .m_peripheral_ar_size(m_peripheral_ar_size),
    .m_peripheral_ar_burst(m_peripheral_ar_burst),
    .m_peripheral_ar_lock(m_peripheral_ar_lock),
    .m_peripheral_ar_cache(m_peripheral_ar_cache),
    .m_peripheral_ar_prot(m_peripheral_ar_prot),
    .m_peripheral_ar_qos(m_peripheral_ar_qos),
    .m_peripheral_r_ready(m_peripheral_r_ready),
    .m_peripheral_r_valid(m_peripheral_r_valid),
    .m_peripheral_r_id(m_peripheral_r_id),
    .m_peripheral_r_data(m_peripheral_r_data),
    .m_peripheral_r_resp(m_peripheral_r_resp),
    .m_peripheral_r_last(m_peripheral_r_last),
    .m_memory_aw_ready(m_memory_aw_ready),
    .m_memory_aw_valid(m_memory_aw_valid),
    .m_memory_aw_id(m_memory_aw_id),
    .m_memory_aw_addr(m_memory_aw_addr),
    .m_memory_aw_len(m_memory_aw_len),
    .m_memory_aw_size(m_memory_aw_size),
    .m_memory_aw_burst(m_memory_aw_burst),
    .m_memory_aw_lock(m_memory_aw_lock),
    .m_memory_aw_cache(m_memory_aw_cache),
    .m_memory_aw_prot(m_memory_aw_prot),
    .m_memory_aw_qos(m_memory_aw_qos),
    .m_memory_w_ready(m_memory_w_ready),
    .m_memory_w_valid(m_memory_w_valid),
    .m_memory_w_data(m_memory_w_data),
    .m_memory_w_strb(m_memory_w_strb),
    .m_memory_w_last(m_memory_w_last),
    .m_memory_b_ready(m_memory_b_ready),
    .m_memory_b_valid(m_memory_b_valid),
    .m_memory_b_id(m_memory_b_id),
    .m_memory_b_resp(m_memory_b_resp),
    .m_memory_ar_ready(m_memory_ar_ready),
    .m_memory_ar_valid(m_memory_ar_valid),
    .m_memory_ar_id(m_memory_ar_id),
    .m_memory_ar_addr(m_memory_ar_addr),
    .m_memory_ar_len(m_memory_ar_len),
    .m_memory_ar_size(m_memory_ar_size),
    .m_memory_ar_burst(m_memory_ar_burst),
    .m_memory_ar_lock(m_memory_ar_lock),
    .m_memory_ar_cache(m_memory_ar_cache),
    .m_memory_ar_prot(m_memory_ar_prot),
    .m_memory_ar_qos(m_memory_ar_qos),
    .m_memory_r_ready(m_memory_r_ready),
    .m_memory_r_valid(m_memory_r_valid),
    .m_memory_r_id(m_memory_r_id),
    .m_memory_r_data(m_memory_r_data),
    .m_memory_r_resp(m_memory_r_resp),
    .m_memory_r_last(m_memory_r_last),
    .io_clock(io_clock),
    .io_reset(io_reset),
    .io_extIntrs(io_extIntrs),
    .io_systemjtag_jtag_TCK(io_systemjtag_jtag_TCK),
    .io_systemjtag_jtag_TMS(io_systemjtag_jtag_TMS),
    .io_systemjtag_jtag_TDI(io_systemjtag_jtag_TDI),
    .io_systemjtag_jtag_TDO_data(io_systemjtag_jtag_TDO_data),
    .io_systemjtag_jtag_TDO_driven(io_systemjtag_jtag_TDO_driven),
    .io_systemjtag_reset(io_systemjtag_reset),
    .io_systemjtag_mfr_id(io_systemjtag_mfr_id),
    .io_systemjtag_part_number(io_systemjtag_part_number),
    .io_systemjtag_version(io_systemjtag_version),
    .io_debug_reset(io_debug_reset),
    .io_riscv_halt_0(io_riscv_halt_0),
    .io_riscv_halt_1(io_riscv_halt_1),
    .scan_mode(scan_mode),
    .dft_lgc_rst_n(dft_lgc_rst_n),
    .dft_mode(dft_mode),
    .dft_ram_hold(dft_ram_hold),
    .dft_ram_bypass(dft_ram_bypass),
    .dft_ram_bp_clken(dft_ram_bp_clken),
    .dft_l3dataram_clk(dft_l3dataram_clk),
    .dft_l3dataramclk_bypass(dft_l3dataramclk_bypass),
    .dft_cgen(dft_cgen)
);
  `include "mem_conn.v"

  tl_monitor_collect#(.SIZE_WD(3),.ADDR_WD(36),.DATA_WD(256),
  .SOURCE_WD(9),.SINK_WD(6),.USER_WD(8),.ECHO_WD(8)
  )tl_monitor_set(
    .clock(io_clock)
  );
endmodule